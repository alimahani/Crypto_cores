`timescale 1ns / 1ps
// ----------------------------------------------------------------------
// Copyright 
// 
// 
//
// ----------------------------------------------------------------------
//----------------------------------------------------------------------------
// Filename:			aes_shiftrow.sv
// Version:				1.00
// Description:	
//
//
// Author:              A. MAHANI
// History:				
//-----------------------------------------------------------------------------

module aes_shiftrow(
                    input    logic [127:0] di,
	                output   logic [127:0] do1);

wire [31:0] r0,r1,r2,r3;
wire [31:0] c0,c1,c2,c3;    
		    
//the original state matrix
//	wire [31:0] r0 = {di[7:0], di[39:32], di[71:64], di[103:96]};
//	wire [31:0] r1 = {di[15:8], di[47:40], di[79:72], di[111, 104]}; 
//	wire [31:0] r2 = {di[23:16], di[55:48], di[87:80], di[119:112]};
//	wire [31:0] r3 = {di[31:24], di[63:56], di[95:88], di[127:120]};

//the state matrix after shift row
assign r0 = {di[7:0],     di[39:32],   di[71:64],   di[103:96]};
assign r1 = {di[47:40],   di[79:72],   di[111:104], di[15:8]  }; 
assign r2 = {di[87:80],   di[119:112], di[23:16],   di[55:48] };
assign r3 = {di[127:120], di[31:24],   di[63:56],   di[95:88] };



assign c0 = {r3[7:0],   r2[7:0],   r1[7:0],   r0[7:0]};
assign c1 = {r3[15:8],  r2[15:8],  r1[15:8],  r0[15:8]};
assign c2 = {r3[23:16], r2[23:16], r1[23:16], r0[23:16]};
assign c3 = {r3[31:24], r2[31:24], r1[31:24], r0[31:24]};
	
	assign do1 = {c3, c0, c1, c2};
	
endmodule