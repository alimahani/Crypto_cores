`timescale 1ns / 1ps
// ----------------------------------------------------------------------
// Copyright 
// 
// 
//
// ----------------------------------------------------------------------
//----------------------------------------------------------------------------
// Filename:			gf_mul3.sv
// Version:				1.00
// Description:	
//
//
// Author:              A. MAHANI
// History:				
//-----------------------------------------------------------------------------

module gf_mul3 (
       input  logic [7:0] di,
       output logic [7:0] do1 );


   logic [7:0] 	      mul2;


   gf_mul2 gf_mul2_0 (.di(di),
	      .do1(mul2));

 
   assign do1 = mul2 ^ di;

endmodule